* c:\users\kumar\esim-workspace\dickson_ckt\dickson_ckt.cir

.lib "sky130_fd_pr/models/sky130.lib.spice" tt


xm1 in in v1 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm2 v1 v1 v2 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm3 v2 v2 v3 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm4 v3 v3 v4 gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xm5 v4 v4 out gnd sky130_fd_pr__nfet_01v8 w=1 l=0.18
xc1  v1 clk1 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xc2  v2 clk2 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xc3  v3 clk1 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xc4  v4 clk2 sky130_fd_pr__cap_mim_m3_1 w=1 l=100
xcout1  out gnd sky130_fd_pr__cap_mim_m3_1 w=1 l=100
v2  clk1 gnd pulse(0 1.8 10n 0 0 10n 20n)
v3  clk2 gnd pulse(0 1.8 0 0 0 10n 20n)
v1 in gnd  dc 1.8
xr1  out gnd gnd sky130_fd_pr__res_high_po_0p69 l=100000
* u1  out plot_v1
.tran 1e-09 100000e-09 0e-00

* Control Statements 
.control
run
print allv > plot_data_v.txt
print alli > plot_data_i.txt
plot v(out)
.endc
.end
